//-------------------------------------------------------------------------------------------------
module dpr
//-------------------------------------------------------------------------------------------------
#
(
	parameter DW = 8,
	parameter AW = 14
)
(
	input  wire         clock1,
	input  wire         ce1,
	output reg [   7:0] q1,
	input  wire[AW-1:0] a1,
	input  wire         clock2,
	input  wire         ce2,
	input  wire         we2,
	input  wire[   7:0] d2,
	output reg [   7:0] q2,
	input  wire[AW-1:0] a2
);
//-------------------------------------------------------------------------------------------------

reg[7:0] d[(2**AW)-1:0];

always @(posedge clock1) if(ce1) q1 <= d[a1];
always @(posedge clock2) if(ce2) if(!we2) d[a2] <= d2; else q2 <= d[a2];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
