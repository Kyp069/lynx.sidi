//-------------------------------------------------------------------------------------------------
module audio
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      reset,
	input  wire      ear,
	input  wire[5:0] dac,
	output wire[1:0] audio
);
//-------------------------------------------------------------------------------------------------

reg source;
always @(posedge clock) source <= ~source;

wire[5:0] mix = source ? {6{ear}} : dac;

//-------------------------------------------------------------------------------------------------

wire q;

dac #(.MSBI(5)) Dac
(
	.clock(clock  ),
	.reset(reset  ),
	.d    (mix    ),
	.q    (q      )
);

assign audio = {2{q}};

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
